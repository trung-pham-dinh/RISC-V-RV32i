`ifndef SINGLECYCLE_SVH
`define SINGLECYCLE_SVH

// `define INST_MEM_PATH "./../02_test/dump/all_inst_and_lsu.mem"
// `define INST_MEM_PATH "./../02_test/dump/stopwatch.mem"
// `define INST_MEM_PATH "./../02_test/dump/all_alu.mem"
// `define INST_MEM_PATH "./../02_test/dump/datmem.mem"
`define INST_MEM_PATH "./../02_test/dump/distance.mem"

`endif
